-- ! comment